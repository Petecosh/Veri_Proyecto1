class scoreboard();
    
endclass