class checkr #(parameter devices = 4);
    pck_drv_chkr paquete_chkr[devices];
    tipo_mbx_drv_chkr drv_chkr_mbx[devices];



endclass