class checker_c;

endclass